module uart_mcu_slavefifo(
    input  sys_clk  ,
    input  sys_rst_n,
    
    input  uart_rxd,
    output uart_txd,

    inout [7:0] cy_D,
    inout [7:0] cy_B,
    input cy_SCL,
    input cy_SDA,
    //input cy_IFCLK                     ,
    //input cy_to_fpga_CTL0_FLAGA        ,
    //input cy_to_fpga_CTL2_FLAGC        ,
    //input cy_to_fpga_CTL1_FLAGB        ,
    //input cy_to_fpga_A7_FLAGD          ,
    output reg cy_from_fpga_RDY1_SLWR       ,//output
    output reg cy_from_fpga_RDY0_SLRD       ,//output
    output reg cy_from_fpga_A2_SLOE         ,//output
    input cy_A0_INT0                   ,// in from pc
    output reg cy_A1_INT1                   ,// out to pc
    input cy_A3_WU2                    ,
    output reg cy_from_fpga_A4_FIFOADR0     ,//output
    output reg cy_from_fpga_A5_FIFOADR1     ,//output
    output reg cy_from_fpga_A6_PKTEND       ,//output

	output reg [7:0] cy_cmd,
	output reg [7:0] cy_dat,
	output reg [7:0] cy_snd_data0,
	output reg [7:0] cy_snd_data1,

    output busy,
    //output [7:0] debug_port0,
    //output [7:0] debug_port1,
    //output [7:0] debug_port2,
    //output debug_pin0,
    //output debug_pin1,
    //output debug_pin2,
    //output debug_pin3,
    //output debug_pin6,
    //output debug_pin7,

    /*
  .sdram_clk_out     (sdram_clk_out),
  .sdram_cke			(sdram_cke),		//SDRAM 时钟有效
  .sdram_cs_n			(sdram_cs_n),		//SDRAM 片选
  .sdram_ras_n		(sdram_ras_n),		//SDRAM 行有效	
  .sdram_cas_n		(sdram_cas_n),		//SDRAM 列有效
  .sdram_we_n			(sdram_we_n),		//SDRAM 写有效
  .sdram_ba			  (sdram_ba),			//SDRAM Bank地址
  .sdram_addr			(sdram_addr),		//SDRAM 行/列地址
  .sdram_data			(sdram_data),		//SDRAM 数据	
  .sdram_dqm		(sdram_dqm),
  .sdram_prob_refresh (sdram_prob_refresh),
*/
    
    //SDRAM 芯片接口
    output        sdram_clk_out,            //SDRAM 芯片时钟
    output        sdram_cke,                //SDRAM 时钟有效
    output        sdram_cs_n,               //SDRAM 片选
    output        sdram_ras_n,              //SDRAM 行有效
    output        sdram_cas_n,              //SDRAM 列有效
    output        sdram_we_n,               //SDRAM 写有效
    output [ 1:0] sdram_ba,                 //SDRAM Bank地址
    output [12:0] sdram_addr,               //SDRAM 行/列地址
    inout  [15:0] sdram_data,               //SDRAM 数据
    output [ 1:0] sdram_dqm,                //SDRAM 数据掩码

    //SDRAM2m 芯片接口
    output        sdram2m_clk_out,            //SDRAM 芯片时钟
    output        sdram2m_cke,                //SDRAM 时钟有效
    output        sdram2m_cs_n,               //SDRAM 片选
    output        sdram2m_ras_n,              //SDRAM 行有效
    output        sdram2m_cas_n,              //SDRAM 列有效
    output        sdram2m_we_n,               //SDRAM 写有效
    output        sdram2m_ba,                 //SDRAM Bank地址
    output [10:0] sdram2m_addr,               //SDRAM 行/列地址
    inout  [15:0] sdram2m_data,               //SDRAM 数据

    
		output reg out_clk,
		output reg out_rst,

		input [7:0] in_pin0,
		input [7:0] in_pin1,
		input [7:0] in_pin2,
		input [7:0] in_pin3,
		input [7:0] in_pin4,
		input [7:0] in_pin5,
		input [7:0] in_pin6,
		input [7:0] in_pin7,

		output reg [7:0] out_pin0,
		output reg [7:0] out_pin1,
		output reg [7:0] out_pin2,
		output reg [7:0] out_pin3,
		output reg [7:0] out_pin4,
		output reg [7:0] out_pin5,
		output reg [7:0] out_pin6,
		output reg [7:0] out_pin7

		);

assign busy = command != 0 && command_done==0;
    
assign cy_D = cy_out_to_pc ? cy_D_out : 8'hzz;
assign cy_B = cy_out_to_pc ? cy_B_out : 8'hzz;
reg [7:0] cy_D_out;
reg [7:0] cy_B_out;

reg cy_out_to_pc;


reg cy_rec_req;
reg cy_snd_ack;
reg [4:0]cy_rec_cnt;
reg [4:0]cy_snd_cnt;
always @(posedge cy_A3_WU2 or negedge sys_rst_n) begin
  if (!sys_rst_n) begin
    cy_cmd<=0;
    cy_dat<=0;
    cy_rec_cnt<=0;
    cy_rec_req<=0;
    cy_snd_ack<=0;
    cy_A1_INT1<=0;
  end else begin
    if         (cy_rec_cnt==0)begin
      if(cy_A0_INT0 && !cy_rec_req)begin
        cy_rec_cnt<=1;
      end
    end else if(cy_rec_cnt==1 )begin cy_cmd[0] <= cy_A0_INT0;cy_rec_cnt<=2;
    end else if(cy_rec_cnt==2 )begin cy_cmd[1] <= cy_A0_INT0;cy_rec_cnt<=3;
    end else if(cy_rec_cnt==3 )begin cy_cmd[2] <= cy_A0_INT0;cy_rec_cnt<=4;
    end else if(cy_rec_cnt==4 )begin cy_cmd[3] <= cy_A0_INT0;cy_rec_cnt<=5;
    end else if(cy_rec_cnt==5 )begin cy_cmd[4] <= cy_A0_INT0;cy_rec_cnt<=6;
    end else if(cy_rec_cnt==6 )begin cy_cmd[5] <= cy_A0_INT0;cy_rec_cnt<=7;
    end else if(cy_rec_cnt==7 )begin cy_cmd[6] <= cy_A0_INT0;cy_rec_cnt<=8;
    end else if(cy_rec_cnt==8 )begin cy_cmd[7] <= cy_A0_INT0;cy_rec_cnt<=9;

    end else if(cy_rec_cnt==9 )begin cy_dat[0] <= cy_A0_INT0;cy_rec_cnt<=10;
    end else if(cy_rec_cnt==10)begin cy_dat[1] <= cy_A0_INT0;cy_rec_cnt<=11;
    end else if(cy_rec_cnt==11)begin cy_dat[2] <= cy_A0_INT0;cy_rec_cnt<=12;
    end else if(cy_rec_cnt==12)begin cy_dat[3] <= cy_A0_INT0;cy_rec_cnt<=13;
    end else if(cy_rec_cnt==13)begin cy_dat[4] <= cy_A0_INT0;cy_rec_cnt<=14;
    end else if(cy_rec_cnt==14)begin cy_dat[5] <= cy_A0_INT0;cy_rec_cnt<=15;
    end else if(cy_rec_cnt==15)begin cy_dat[6] <= cy_A0_INT0;cy_rec_cnt<=16;
    end else if(cy_rec_cnt==16)begin cy_dat[7] <= cy_A0_INT0;cy_rec_cnt<=0;cy_rec_req<=1;
    end

    if(cy_snd_req && !cy_snd_ack)begin
      if         (cy_snd_cnt==0 )begin cy_snd_cnt<=1 ;cy_A1_INT1 <= 1;
      
      end else if(cy_snd_cnt==1 )begin cy_snd_cnt<=2 ;cy_A1_INT1 <= cy_snd_data0[0];
      end else if(cy_snd_cnt==2 )begin cy_snd_cnt<=3 ;cy_A1_INT1 <= cy_snd_data0[1];
      end else if(cy_snd_cnt==3 )begin cy_snd_cnt<=4 ;cy_A1_INT1 <= cy_snd_data0[2];
      end else if(cy_snd_cnt==4 )begin cy_snd_cnt<=5 ;cy_A1_INT1 <= cy_snd_data0[3];
      end else if(cy_snd_cnt==5 )begin cy_snd_cnt<=6 ;cy_A1_INT1 <= cy_snd_data0[4];
      end else if(cy_snd_cnt==6 )begin cy_snd_cnt<=7 ;cy_A1_INT1 <= cy_snd_data0[5];
      end else if(cy_snd_cnt==7 )begin cy_snd_cnt<=8 ;cy_A1_INT1 <= cy_snd_data0[6];
      end else if(cy_snd_cnt==8 )begin cy_snd_cnt<=9 ;cy_A1_INT1 <= cy_snd_data0[7];

      end else if(cy_snd_cnt==9 )begin cy_snd_cnt<=10;cy_A1_INT1 <= cy_snd_data1[0];
      end else if(cy_snd_cnt==10)begin cy_snd_cnt<=11;cy_A1_INT1 <= cy_snd_data1[1];
      end else if(cy_snd_cnt==11)begin cy_snd_cnt<=12;cy_A1_INT1 <= cy_snd_data1[2];
      end else if(cy_snd_cnt==12)begin cy_snd_cnt<=13;cy_A1_INT1 <= cy_snd_data1[3];
      end else if(cy_snd_cnt==13)begin cy_snd_cnt<=14;cy_A1_INT1 <= cy_snd_data1[4];
      end else if(cy_snd_cnt==14)begin cy_snd_cnt<=15;cy_A1_INT1 <= cy_snd_data1[5];
      end else if(cy_snd_cnt==15)begin cy_snd_cnt<=16;cy_A1_INT1 <= cy_snd_data1[6];
      end else if(cy_snd_cnt==16)begin cy_snd_cnt<=17;cy_A1_INT1 <= cy_snd_data1[7];
      end else if(cy_snd_cnt==17)begin cy_snd_cnt<=18;cy_A1_INT1 <= 0;cy_snd_ack<=1;
      end
    end else begin
      cy_snd_cnt<=0;
      cy_snd_ack<=0;
    end

    
    if(cy_rec_req && cy_rec_ack)begin
      cy_rec_req<=0;
    end
    
    
    
  end
end









    
wire uart_rec;
wire [7:0] uart_data_r;
reg uart_send;
reg [7:0] uart_data_w;

reg [7:0] uw_reg0;
reg [7:0] uw_reg1;
reg [7:0] uw_reg2;
reg [7:0] uw_reg3;
reg [7:0] uw_reg4;
reg [7:0] uw_reg5;
reg [7:0] uw_reg6;
reg [7:0] uw_reg7;

reg [7:0] ur_reg0;
reg [7:0] ur_reg1;
reg [7:0] ur_reg2;
reg [7:0] ur_reg3;
reg [7:0] ur_reg4;
reg [7:0] ur_reg5;
reg [7:0] ur_reg6;
reg [7:0] ur_reg7;

reg uart_rec_last;
wire uart_rec_rise;
assign uart_rec_rise = uart_rec && !uart_rec_last;
always @(posedge sys_clk or negedge sys_rst_n) begin
  if (!sys_rst_n) begin
		uart_rec_last<=0;
  end else begin
		uart_rec_last <= uart_rec;
	end
end
///////////
uart_hs ins_uart_hs(
    .sys_clk        (sys_clk), 
    .sys_rst_n      (sys_rst_n),
    .uart_rxd       (uart_rxd),
    .uart_txd       (uart_txd),

    .uart_rec       (uart_rec),
    .uart_data_out  (uart_data_r),
    .uart_send      (uart_send),
    .uart_data_in   (uart_data_w)
  );

  
reg cy_rec_ack;
reg [7:0] command;
reg [7:0] data;
reg [15:0] data_index;
reg data_arrive;
reg cy_rec_req_buff;
always @(posedge sys_clk or negedge sys_rst_n) begin
  if (!sys_rst_n) begin
    command <= 0;
    data <= 0;
    data_index<=0;
    data_arrive<=0;
    cy_rec_ack<=0;
  end else begin
	cy_rec_req_buff<=cy_rec_req;
    data_arrive <= 0;
    if (uart_rec_rise) begin //串口数据到达
      if(command==8'b0) begin
        command <= uart_data_r;
        data_index <= 16'hFFFF;
      end else begin
        data_arrive <= 1;
        data_index <= data_index + 1'b1;
        data <= uart_data_r;
      end
    end
    
    if(!cy_rec_req_buff && cy_rec_ack)begin
      cy_rec_ack <= 0;
    end
    
    if (cy_rec_req_buff && !cy_rec_ack) begin //cy数据到达
      command <= cy_cmd;
      cy_rec_ack <= 1;
    end
    if(command_done)begin
      command <= 0;
    end
  end
end

reg command_done;
reg [10:0] timer;
reg [7:0] reg_temp;
reg [9:0] timer2;
reg [23:0] read_address;
reg hibit;

reg [15:0] timer3;

reg [7:0] sum;
reg [15:0] sum16;

reg cy_snd_req;

reg [16:0] temp_val;
always @(posedge sys_clk or negedge sys_rst_n) begin
  if (!sys_rst_n) begin
    out_pin0<=8'bzzzzzzzz;
    out_pin1<=8'bzzzzzzzz;
    out_pin2<=8'bzzzzzzzz;
    out_pin3<=8'bzzzzzzzz;
    out_pin4<=8'bzzzzzzzz;
    out_pin5<=8'bzzzzzzzz;
    out_pin6<=8'bzzzzzzzz;
    out_pin7<=8'bzzzzzzzz;
    
    uw_reg0<=0;
    uw_reg1<=0;
    uw_reg2<=0;
    uw_reg3<=0;
    uw_reg4<=0;
    uw_reg5<=0;
    uw_reg6<=0;
    uw_reg7<=0;
    
    uart_send<=0;
    uart_data_w<=0;
    out_clk<=0;
    out_rst<=0;
    command_done <= 0;
    timer<=0;
    timer2<=0;
    timer3<=0;
    sdram_c_address <= 0;
    sdram_c_data_in <= 0;
    sdram_c_read_req <= 0;
    sdram_c_write_req <= 0;
    sdram_c_write_en <= 0;
    sdram_c_write_latch_address <=0;
    sum <=0;
	 sum16 <=0;


    cy_from_fpga_A2_SLOE<=1;
    cy_from_fpga_RDY0_SLRD<=1;
    cy_from_fpga_RDY1_SLWR<=1;
    cy_from_fpga_A4_FIFOADR0<=0;
    cy_from_fpga_A5_FIFOADR1<=0;
    cy_from_fpga_A6_PKTEND<=1;
		
	 cy_out_to_pc<=0;
	
    cy_snd_req<=0;
    cy_snd_data0 <= 0;
    cy_snd_data1 <= 0;

  end else begin

    if(cy_snd_ack)begin
      cy_snd_req <= 0;
    end
    
    if(command_done)begin
      uart_send<=0;
      if          (command == 8'h00) begin 
        command_done<=0;
      end
    end else begin//command_done==0
      if          (command == 8'h00) begin
      end else if (command == 8'h10) begin out_clk<=1; command_done<=1;
      end else if (command == 8'h11) begin out_clk<=0; command_done<=1;
      end else if (command == 8'h12) begin out_rst<=1; command_done<=1;
      end else if (command == 8'h13) begin out_rst<=0; command_done<=1;

      end else if (command == 8'h20) begin uart_send<=1; uart_data_w<=in_pin0; command_done<=1;
      end else if (command == 8'h21) begin uart_send<=1; uart_data_w<=in_pin1; command_done<=1;
      end else if (command == 8'h22) begin uart_send<=1; uart_data_w<=in_pin2; command_done<=1;
      end else if (command == 8'h23) begin uart_send<=1; uart_data_w<=in_pin3; command_done<=1;
      end else if (command == 8'h24) begin uart_send<=1; uart_data_w<=in_pin4; command_done<=1;
      end else if (command == 8'h25) begin uart_send<=1; uart_data_w<=in_pin5; command_done<=1;
      end else if (command == 8'h26) begin uart_send<=1; uart_data_w<=in_pin6; command_done<=1;
      end else if (command == 8'h27) begin uart_send<=1; uart_data_w<=in_pin7; command_done<=1;

      end else if (command == 8'h30) begin if(data_arrive)begin out_pin0<=data; command_done<=1;end
      end else if (command == 8'h31) begin if(data_arrive)begin out_pin1<=data; command_done<=1;end
      end else if (command == 8'h32) begin if(data_arrive)begin out_pin2<=data; command_done<=1;end
      end else if (command == 8'h33) begin if(data_arrive)begin out_pin3<=data; command_done<=1;end
      end else if (command == 8'h34) begin if(data_arrive)begin out_pin4<=data; command_done<=1;end
      end else if (command == 8'h35) begin if(data_arrive)begin out_pin5<=data; command_done<=1;end
      end else if (command == 8'h36) begin if(data_arrive)begin out_pin6<=data; command_done<=1;end
      end else if (command == 8'h37) begin if(data_arrive)begin out_pin7<=data; command_done<=1;end

      end else if (command == 8'h40) begin if(data_arrive)begin uw_reg0<=data; command_done<=1;end
      end else if (command == 8'h41) begin if(data_arrive)begin uw_reg1<=data; command_done<=1;end
      end else if (command == 8'h42) begin if(data_arrive)begin uw_reg2<=data; command_done<=1;end
      end else if (command == 8'h43) begin if(data_arrive)begin uw_reg3<=data; command_done<=1;end
      end else if (command == 8'h44) begin if(data_arrive)begin uw_reg4<=data; command_done<=1;end
      end else if (command == 8'h45) begin if(data_arrive)begin uw_reg5<=data; command_done<=1;end
      end else if (command == 8'h46) begin if(data_arrive)begin uw_reg6<=data; command_done<=1;end
      end else if (command == 8'h47) begin if(data_arrive)begin uw_reg7<=data; command_done<=1;end

      end else if (command == 8'h50) begin uart_send<=1; uart_data_w<=ur_reg0; command_done<=1;
      end else if (command == 8'h51) begin uart_send<=1; uart_data_w<=ur_reg1; command_done<=1;
      end else if (command == 8'h52) begin uart_send<=1; uart_data_w<=ur_reg2; command_done<=1;
      end else if (command == 8'h53) begin uart_send<=1; uart_data_w<=ur_reg3; command_done<=1;
      end else if (command == 8'h54) begin uart_send<=1; uart_data_w<=ur_reg4; command_done<=1;
      end else if (command == 8'h55) begin uart_send<=1; uart_data_w<=ur_reg5; command_done<=1;
      end else if (command == 8'h56) begin uart_send<=1; uart_data_w<=ur_reg6; command_done<=1;
      end else if (command == 8'h57) begin uart_send<=1; uart_data_w<=ur_reg7; command_done<=1;

      end else if (command == 8'h60) begin out_pin0<=8'bzzzzzzzz; command_done<=1;
      end else if (command == 8'h61) begin out_pin1<=8'bzzzzzzzz; command_done<=1;
      end else if (command == 8'h62) begin out_pin2<=8'bzzzzzzzz; command_done<=1;
      end else if (command == 8'h63) begin out_pin3<=8'bzzzzzzzz; command_done<=1;
      end else if (command == 8'h64) begin out_pin4<=8'bzzzzzzzz; command_done<=1;
      end else if (command == 8'h65) begin out_pin5<=8'bzzzzzzzz; command_done<=1;
      end else if (command == 8'h66) begin out_pin6<=8'bzzzzzzzz; command_done<=1;
      end else if (command == 8'h67) begin out_pin7<=8'bzzzzzzzz; command_done<=1;

      end else if (command == 8'h70) begin uw_reg0<=cy_dat; command_done<=1;
      end else if (command == 8'h71) begin uw_reg1<=cy_dat; command_done<=1;
      end else if (command == 8'h72) begin uw_reg2<=cy_dat; command_done<=1;
      end else if (command == 8'h73) begin uw_reg3<=cy_dat; command_done<=1;
      end else if (command == 8'h74) begin uw_reg4<=cy_dat; command_done<=1;
      end else if (command == 8'h75) begin uw_reg5<=cy_dat; command_done<=1;
      end else if (command == 8'h76) begin uw_reg6<=cy_dat; command_done<=1;
      end else if (command == 8'h77) begin uw_reg7<=cy_dat; command_done<=1;

      end else if (command == 8'hA0) begin//sdram write
        timer<=timer+1'b1;
        if(timer==0)begin
          sdram_c_address <= {uw_reg4,uw_reg3,uw_reg2};
          sdram_c_data_in <= {uw_reg1,uw_reg0};
          sdram_c_write_req<=1;
        end else begin
          if(sdram_c_write_ack)begin
            ur_reg7<=timer[7:0];
            timer<=0;
            sdram_c_write_req<=0;
            command_done<=1;
          end
        end

      end else if (command == 8'hA1) begin//sdram read
        timer<=timer+1'b1;
        if(timer==0)begin
          sdram_c_address <= {uw_reg4,uw_reg3,uw_reg2};
          sdram_c_read_req<=1;
        end else begin
          if(sdram_c_read_ack)begin
            ur_reg7 <= timer[7:0];
            timer <= 0;
            ur_reg0 <= sdram_c_data_out[7:0];
            ur_reg1 <= sdram_c_data_out[15:8];
            sdram_c_read_req<=0;
            command_done <= 1;
          end
        end

      end else if (command == 8'hA2) begin//sdram long write
        if(data_arrive)begin
          if (data_index[0]==0)begin
            reg_temp <= data;//锁存低字节
          end else begin
            sdram_c_write_en <= 1;
            sdram_c_data_in<={data,reg_temp};
            if         (data_index==1)begin
              sdram_c_write_latch_address <= 1;
              sdram_c_address <= {uw_reg4,uw_reg3,uw_reg2};
            end else if(data_index==513)begin
              sdram_c_write_en <= 0;
              uart_send<=1;
              uart_data_w<=8'h41;//'A' 8'h41;
              command_done <= 1;
            end
          end
        end else begin
          sdram_c_write_en <= 0;
          sdram_c_write_latch_address <= 0;
        end

      end else if (command == 8'hA3) begin//sdram long read
        timer2<=timer2+1'b1;
        uart_send<=0;
        if(timer2==600)begin//25 * 10 +50
          timer2<=0;
        end
        if(timer2==0)begin
          if(timer==0)begin//锁存地址
            read_address    <= {uw_reg4,uw_reg3,uw_reg2};
            sdram_c_address <= {uw_reg4,uw_reg3,uw_reg2};
            sum <= 0;
          end else begin
            if(timer[0]==1)begin
              read_address <= read_address+1'b1;
            end
            sdram_c_address <= read_address;
          end
          sdram_c_read_req<=1;
        end else begin
          if(sdram_c_read_req && sdram_c_read_ack)begin
            timer<=timer+1'b1;
            sdram_c_read_req<=0;
            sum <= sum + ((timer[0]==1)?sdram_c_data_out[15:8]:sdram_c_data_out[7:0]);
            uart_send<=1;
            uart_data_w<=(timer[0]==1)?sdram_c_data_out[15:8]:sdram_c_data_out[7:0];
            if(timer==1024)begin
              uart_send<=1;
              uart_data_w<=sum;
              timer2<=0;
              timer<=0;
              command_done<=1;
            end
          end
        end
        
 
      end else if (command == 8'hB0) begin//sdram long write ok
        timer3 <= timer3 + 1'b1;
        sdram_c_write_latch_address<=0;

        if         (timer3==0)begin																	//step0
          cy_from_fpga_A2_SLOE<=0;//on
          cy_from_fpga_RDY0_SLRD<=0;//on
          sdram_c_address <= {uw_reg4,uw_reg3,uw_reg2};
        end else if(timer3==(512 * 4 + 2))begin																	//step5  n字*4+2
          cy_from_fpga_A2_SLOE<=1;//off
          cy_from_fpga_RDY0_SLRD<=1;//off
          timer3<=0;
          command_done<=1;
          cy_snd_req <= 1;
          cy_snd_data0 <= 8'h12;
          cy_snd_data1 <= 8'h34;
        end else begin
          if         (timer3[1:0]==1)begin																	//step1
            cy_from_fpga_RDY0_SLRD<=0;//on
          end else if(timer3[1:0]==2)begin																	//step2
            cy_from_fpga_RDY0_SLRD<=1;//off
            //读取 并写入sdram
            sdram_c_write_en<=1;
            if(timer3==2)begin sdram_c_write_latch_address<=1; end
            sdram_c_data_in<={cy_D,cy_B};
          end else if(timer3[1:0]==3)begin																	//step3
            cy_from_fpga_RDY0_SLRD<=1;//off
            sdram_c_write_en<=0;
          end else begin																			//step4
            cy_from_fpga_RDY0_SLRD<=0;//on
            sdram_c_write_en<=0;
          end
        end
        

      end else if (command == 8'hB1) begin//sdram long read
        timer2<=timer2+1'b1;
        
        if(timer2==0)begin
          if(timer==0)begin//锁存地址
            sdram_c_address <= {uw_reg4,uw_reg3,uw_reg2};
            sum16 <= 0;
            cy_from_fpga_A4_FIFOADR0<=0;//set channel
            cy_from_fpga_A5_FIFOADR1<=1;
            cy_out_to_pc<=1;//set out
          end else begin
            sdram_c_address <= sdram_c_address + 1'b1;
            
          end
          sdram_c_read_req<=1;
        end else if(timer2==30) begin//sdram 响应
          if(!sdram_c_read_ack)begin
            //err
          end
          timer<=timer+1'b1;
          sdram_c_read_req<=0;
          sum16 <= sum16 + sdram_c_data_out;
          cy_D_out = sdram_c_data_out[15:8];
          cy_B_out = sdram_c_data_out[7:0];
          cy_from_fpga_RDY1_SLWR<=0;//set wr
 
        end else if(timer2==60)begin
			cy_from_fpga_RDY1_SLWR<=1;//set wr
          if(timer==513)begin
            cy_from_fpga_A4_FIFOADR0<=0;//set channel
            cy_from_fpga_A5_FIFOADR1<=0;
            cy_out_to_pc<=0;//set out
            timer<=0;
            command_done<=1;
            cy_snd_req <= 1;
            cy_snd_data1 <= sum16[15:8];
            cy_snd_data0 <= sum16[7:0];
          end
          timer2<=0;
        end
        
		  

      end else if (command == 8'hC0) begin//sdram2m long write ok
        timer3 <= timer3 + 1'b1;
        sdram2m_c_write_latch_address<=0;

        if         (timer3==0)begin																	//step0
          cy_from_fpga_A2_SLOE<=0;//on
          cy_from_fpga_RDY0_SLRD<=0;//on
          sdram2m_c_address <= {uw_reg4,uw_reg3,uw_reg2};
        end else if(timer3==(512 * 4 + 2))begin																	//step5  n字*4+2
          cy_from_fpga_A2_SLOE<=1;//off
          cy_from_fpga_RDY0_SLRD<=1;//off
          timer3<=0;
          command_done<=1;
          cy_snd_req <= 1;
          cy_snd_data0 <= 8'h12;
          cy_snd_data1 <= 8'h34;
        end else begin
          if         (timer3[1:0]==1)begin																	//step1
            cy_from_fpga_RDY0_SLRD<=0;//on
          end else if(timer3[1:0]==2)begin																	//step2
            cy_from_fpga_RDY0_SLRD<=1;//off
            //读取 并写入sdram2m
            sdram2m_c_write_en<=1;
            if(timer3==2)begin sdram2m_c_write_latch_address<=1; end
            sdram2m_c_data_in<={cy_D,cy_B};
          end else if(timer3[1:0]==3)begin																	//step3
            cy_from_fpga_RDY0_SLRD<=1;//off
            sdram2m_c_write_en<=0;
          end else begin																			//step4
            cy_from_fpga_RDY0_SLRD<=0;//on
            sdram2m_c_write_en<=0;
          end
        end
        

      end else if (command == 8'hC1) begin//sdram2m long read
        timer2<=timer2+1'b1;
        
        if(timer2==0)begin
          if(timer==0)begin//锁存地址
            sdram2m_c_address <= {uw_reg4,uw_reg3,uw_reg2};
            sum16 <= 0;
            cy_from_fpga_A4_FIFOADR0<=0;//set channel
            cy_from_fpga_A5_FIFOADR1<=1;
            cy_out_to_pc<=1;//set out
          end else begin
            sdram2m_c_address <= sdram2m_c_address + 1'b1;
            
          end
          sdram2m_c_read_req<=1;
        end else if(timer2==30) begin//sdram2m 响应
          if(!sdram2m_c_read_ack)begin
            //err
          end
          timer<=timer+1'b1;
          sdram2m_c_read_req<=0;
          sum16 <= sum16 + sdram2m_c_data_out;
          cy_D_out = sdram2m_c_data_out[15:8];
          cy_B_out = sdram2m_c_data_out[7:0];
          cy_from_fpga_RDY1_SLWR<=0;//set wr
 
        end else if(timer2==60)begin
			cy_from_fpga_RDY1_SLWR<=1;//set wr
          if(timer==513)begin
            cy_from_fpga_A4_FIFOADR0<=0;//set channel
            cy_from_fpga_A5_FIFOADR1<=0;
            cy_out_to_pc<=0;//set out
            timer<=0;
            command_done<=1;
            cy_snd_req <= 1;
            cy_snd_data1 <= sum16[15:8];
            cy_snd_data0 <= sum16[7:0];
          end
          timer2<=0;
        end
                
        
      end
    end
  end
end









reg [23:0] sdram_c_address;
reg [15:0] sdram_c_data_in;
wire [15:0] sdram_c_data_out;
reg  sdram_c_read_req;
wire  sdram_c_read_ack;
reg  sdram_c_write_req;
wire  sdram_c_write_ack;
reg sdram_c_write_en;
reg sdram_c_write_latch_address;
sdram ins_sdram(
  .sys_clk    (sys_clk  ),       // 时钟信号
  .sys_rst_n  (sys_rst_n),       // 复位信号

  //SDRAM 芯片接口
  .sdram_clk_out     (sdram_clk_out),
  .sdram_cke			(sdram_cke),		//SDRAM 时钟有效
  .sdram_cs_n			(sdram_cs_n),		//SDRAM 片选
  .sdram_ras_n		(sdram_ras_n),		//SDRAM 行有效	
  .sdram_cas_n		(sdram_cas_n),		//SDRAM 列有效
  .sdram_we_n			(sdram_we_n),		//SDRAM 写有效
  .sdram_ba			  (sdram_ba),			//SDRAM Bank地址
  .sdram_addr			(sdram_addr),		//SDRAM 行/列地址
  .sdram_data			(sdram_data),		//SDRAM 数据	
  .sdram_dqm		(sdram_dqm),

  .clk        (sys_clk),//in
  .address    (sdram_c_address),//in
  .data_in    (sdram_c_data_in),//in
  .data_out   (sdram_c_data_out),//out
  .read_req   (sdram_c_read_req),//in
  .read_ack   (sdram_c_read_ack),//out
  .write_req  (sdram_c_write_req),//in
  .write_ack  (sdram_c_write_ack),//out
  .write_en   (sdram_c_write_en),//in
  .write_latch_address(sdram_c_write_latch_address)//in
);


reg [19:0] sdram2m_c_address;
reg [15:0] sdram2m_c_data_in;
wire [15:0] sdram2m_c_data_out;
reg  sdram2m_c_read_req;
wire  sdram2m_c_read_ack;
reg  sdram2m_c_write_req;
wire  sdram2m_c_write_ack;
reg sdram2m_c_write_en;
reg sdram2m_c_write_latch_address;
sdram2m(
  .sys_clk    (sys_clk  ),       // 时钟信号
  .sys_rst_n  (sys_rst_n),       // 复位信号

  //SDRAM 芯片接口
  .sdram_clk_out     (sdram2m_clk_out),
  .sdram_cke			(sdram2m_cke),		//SDRAM 时钟有效
  .sdram_cs_n			(sdram2m_cs_n),		//SDRAM 片选
  .sdram_ras_n		(sdram2m_ras_n),		//SDRAM 行有效	
  .sdram_cas_n		(sdram2m_cas_n),		//SDRAM 列有效
  .sdram_we_n			(sdram2m_we_n),		//SDRAM 写有效
  .sdram_ba			  (sdram2m_ba),			//SDRAM Bank地址
  .sdram_addr			(sdram2m_addr),		//SDRAM 行/列地址
  .sdram_data			(sdram2m_data),		//SDRAM 数据	

  .clk        (sys_clk),//in
  .address    (sdram2m_c_address),//in
  .data_in    (sdram2m_c_data_in),//in
  .data_out   (sdram2m_c_data_out),//out
  .read_req   (sdram2m_c_read_req),//in
  .read_ack   (sdram2m_c_read_ack),//out
  .write_req  (sdram2m_c_write_req),//in
  .write_ack  (sdram2m_c_write_ack),//out
  .write_en   (sdram2m_c_write_en),//in
  .write_latch_address(sdram2m_c_write_latch_address)//in

);


endmodule
